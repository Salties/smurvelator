module stimulus;
initial
begin
    $display("hello,world");
    $finish;
end
endmodule
