module our;
initial
begin
    $display("hello,world");
    $finish;
end
endmodule
